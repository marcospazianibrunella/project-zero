`define DEBUG

`define AXIS_ETH_DATA_WIDTH 512
`define AXIS_ETH_KEEP_WIDTH `AXIS_ETH_DATA_WIDTH / 8
`define AXIS_ETH_SYNC_DATA_WIDTH `AXIS_ETH_DATA_WIDTH
`define AXIS_ETH_TX_USER_WIDTH 1
`define AXIS_ETH_RX_USER_WIDTH 1
